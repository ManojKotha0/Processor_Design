
module Data_Memory 
(
    //input clk,            
    input MemRead,             
    input MemWrite,            
    input [63:0] address,    
    input [63:0] write_data,  
    output reg [63:0] read_data  
);

    reg [63:0] memory [0:255];  
    initial begin
        // memory[0]=64'h0000000000000000;
        // memory[1]=64'h0000000000000001;
        // memory[2]=64'h0000000000000002;
        // memory[3]=64'h0000000000000003;
        // memory[4]=64'h0000000000000004;
        // memory[5]=64'h0000000000000005;
        // memory[6]=64'h0000000000000006;
        // memory[7]=64'h0000000000000007;
        // memory[8]=64'h0000000000000008;
        memory[0]  = 64'h0000000000000000;
        memory[1]  = 64'h0000000000000000;
        memory[2]  = 64'h0000000000000000;
        memory[3]  = 64'h0000000000000000;
        memory[4]  = 64'h0000000000000000;
        memory[5]  = 64'h0000000000000000;
        memory[6]  = 64'h0000000000000000;
        memory[7]  = 64'h0000000000000000;
        memory[8]  = 64'h0000000000000000;
        memory[9]  = 64'h0000000000000000;
        memory[10] = 64'h0000000000000000;
        memory[11] = 64'h0000000000000000;
        memory[12] = 64'h0000000000000000;
        memory[13] = 64'h0000000000000000;
        memory[14] = 64'h0000000000000000;
        memory[15] = 64'h0000000000000000;
        memory[16] = 64'h0000000000000000;
        memory[17] = 64'h0000000000000000;
        memory[18] = 64'h0000000000000000;
        memory[19] = 64'h0000000000000000;
        memory[20] = 64'h0000000000000000;
        memory[21] = 64'h0000000000000000;
        memory[22] = 64'h0000000000000000;
        memory[23] = 64'h0000000000000000;
        memory[24] = 64'h0000000000000000;
        memory[25] = 64'h0000000000000000;
        memory[26] = 64'h0000000000000000;
        memory[27] = 64'h0000000000000000;
        memory[28] = 64'h0000000000000000;
        memory[29] = 64'h0000000000000000;
        memory[30] = 64'h0000000000000000;
        memory[31] = 64'h0000000000000000;
        memory[32] = 64'h0000000000000000;
        memory[33] = 64'h0000000000000000;
        memory[34] = 64'h0000000000000000;
        memory[35] = 64'h0000000000000000;
        memory[36] = 64'h0000000000000000;
        memory[37] = 64'h0000000000000000;
        memory[38] = 64'h0000000000000000;
        memory[39] = 64'h0000000000000000;
        memory[40] = 64'h0000000000000000;
        memory[41] = 64'h0000000000000000;
        memory[42] = 64'h0000000000000000;
        memory[43] = 64'h0000000000000000;
        memory[44] = 64'h0000000000000000;
        memory[45] = 64'h0000000000000000;
        memory[46] = 64'h0000000000000000;
        memory[47] = 64'h0000000000000000;
        memory[48] = 64'h0000000000000000;
        memory[49] = 64'h0000000000000000;
        memory[50] = 64'h0000000000000000;
        memory[51] = 64'h0000000000000000;
        memory[52] = 64'h0000000000000000;
        memory[53] = 64'h0000000000000000;
        memory[54] = 64'h0000000000000000;
        memory[55] = 64'h0000000000000000;
        memory[56] = 64'h0000000000000000;
        memory[57] = 64'h0000000000000000;
        memory[58] = 64'h0000000000000000;
        memory[59] = 64'h0000000000000000;
        memory[60] = 64'h0000000000000000;
        memory[61] = 64'h0000000000000000;
        memory[62] = 64'h0000000000000000;
        memory[63] = 64'h0000000000000000;
        memory[64]  = 64'h0000000000000000;
        memory[65]  = 64'h0000000000000000;
        memory[66]  = 64'h0000000000000000;
        memory[67]  = 64'h0000000000000000;
        memory[68]  = 64'h0000000000000000;
        memory[69]  = 64'h0000000000000000;
        memory[70]  = 64'h0000000000000000;
        memory[71]  = 64'h0000000000000000;
        memory[72]  = 64'h0000000000000000;
        memory[73]  = 64'h0000000000000000;
        memory[74] = 64'h0000000000000000;
        memory[75] = 64'h0000000000000000;
        memory[76] = 64'h0000000000000000;
        memory[77] = 64'h0000000000000000;
        memory[78] = 64'h0000000000000000;
        memory[79] = 64'h0000000000000000;
        memory[80] = 64'h0000000000000000;
        memory[81] = 64'h0000000000000000;
        memory[82] = 64'h0000000000000000;
        memory[83] = 64'h0000000000000000;
        memory[84] = 64'h0000000000000000;
        memory[85] = 64'h0000000000000000;
        memory[86] = 64'h0000000000000000;
        memory[87] = 64'h0000000000000000;
        memory[88] = 64'h0000000000000000;
        memory[89] = 64'h0000000000000000;
        memory[90] = 64'h0000000000000000;
        memory[91] = 64'h0000000000000000;
        memory[92] = 64'h0000000000000000;
        memory[93] = 64'h0000000000000000;
        memory[94] = 64'h0000000000000000;
        memory[95] = 64'h0000000000000000;
        memory[96] = 64'h0000000000000000;
        memory[97] = 64'h0000000000000000;
        memory[98] = 64'h0000000000000000;
        memory[99] = 64'h0000000000000000;
        memory[100] = 64'h0000000000000000;
        memory[101] = 64'h0000000000000000;
        memory[102] = 64'h0000000000000000;
        memory[103] = 64'h0000000000000000;
        memory[104] = 64'h0000000000000000;
        memory[105] = 64'h0000000000000000;
        memory[106] = 64'h0000000000000000;
        memory[107] = 64'h0000000000000000;
        memory[108] = 64'h0000000000000000;
        memory[109] = 64'h0000000000000000;
        memory[110] = 64'h0000000000000000;
        memory[111] = 64'h0000000000000000;
        memory[112] = 64'h0000000000000000;
        memory[113] = 64'h0000000000000000;
        memory[114] = 64'h0000000000000000;
        memory[115] = 64'h0000000000000000;
        memory[116] = 64'h0000000000000000;
        memory[117] = 64'h0000000000000000;
        memory[118] = 64'h0000000000000000;
        memory[119] = 64'h0000000000000000;
        memory[120] = 64'h0000000000000000;
        memory[121] = 64'h0000000000000000;
        memory[122] = 64'h0000000000000000;
        memory[123] = 64'h0000000000000000;
        memory[124] = 64'h0000000000000000;
        memory[125] = 64'h0000000000000000;
        memory[126] = 64'h0000000000000000;
        memory[127] = 64'h0000000000000000;
    end

    
    always @(*) begin
        if (MemWrite) 
            memory[address[9:0]] <= write_data;
        if (MemRead) 
            read_data <= memory[address[9:0]];
    end
    // always @(*) begin
    //     if (MemRead) 
    //         read_data <= memory[address[9:0]];
    // end

endmodule